module rom(
    input wire rst,
    input wire clk,
    input wire [31:0] pc_i,
    
    output reg [31:0] inst_o
);

    reg [31:0] rom[0:3];
    initial $readmemh("E:Documents/bianchengwenjian/mips32-CPU/dev/sources_1/new/rom.data", rom);
    
    always @ (*) begin
        if(rst == 1'b1) begin
            inst_o <= 32'b0;
        end else begin
            inst_o <= rom[pc_i[3:2]];
        end
    end
endmodule

